module ifs #(
    N = 32
) (
    
);
    
endmodule